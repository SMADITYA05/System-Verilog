module func(input int a,b);
  function compare(a,b);
    if(a>b)
      $display("a is greater");
    else if(a==b)
      $display("one and the same");
    else
      $display("b is greater");
  endfunction
  initial begin
    compare(6,9);
    compare(9,6);
    compare(5,5);
  end
endmodule
